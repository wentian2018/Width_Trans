module  width_trans (

    input [3:0] txd_in;
    input tx_en_in;
    input tx_clk_in;//tx_clk_in is 25MHz

    input rstn;

    output [2:0] txd_out;
    output tx_en_out;

    
    input tx_clk_out;//tx_clk_out is 33.3333333...Mhz

);





endmodule


