module  



endmodule


